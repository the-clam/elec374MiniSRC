`timescale 1 ns/10 ps
module alu_div(
	input wire [31:0] A, // divident
   input wire [31:0] B, // divisor
	output wire [31:0] Q
);

endmodule