module 32_to_1_mux(
	// clk
	input clk,
	// registers,
	input [31:0] BusMuxIn_R0,
	input [31:0] BusMuxIn_R1,
	input [31:0] BusMuxIn_R2,
	input [31:0] BusMuxIn_R3,
	input [31:0] BusMuxIn_R4,
	input [31:0] BusMuxIn_R5,
	input [31:0] BusMuxIn_R6,
	input [31:0] BusMuxIn_R7,
	input [31:0] BusMuxIn_R8,
	input [31:0] BusMuxIn_R9,
	input [31:0] BusMuxIn_R10,
	input [31:0] BusMuxIn_R11,
	input [31:0] BusMuxIn_R12,
	input [31:0] BusMuxIn_R13,
	input [31:0] BusMuxIn_R14,
	input [31:0] BusMuxIn_R15,
	// other Inputs
	input [31:0] BusMuxIn_HI,
	input [31:0] BuxMuxIn_LO,
	input [31:0] BuxMuxIn_Zhigh,
	input [31:0] BuxMuxIn_Zlow,
	input [31:0] BuxMuxIn_PC,
	input [31:0] BuxMuxIn_MDR,
	input [31:0] BuxMuxIn_InPort,
	input [31:0] C_sign_extended,

	// mux output
	output [31:0] BusMuxOut,
	
	// Select signal for the multiplexer
	input [4:0] mux_select

);

always@(clk)
begin
	// outputs for each case
	if(mux_select[4:0] == 5'b00000) BusMuxOut[31:0] <= BusMuxIn_R0 [31:0];
	if(mux_select[4:0] == 5'b00001) BusMuxOut[31:0] <= BusMuxIn_R1 [31:0];
	if(mux_select[4:0] == 5'b00010) BusMuxOut[31:0] <= BusMuxIn_R2 [31:0];
	if(mux_select[4:0] == 5'b00011) BusMuxOut[31:0] <= BusMuxIn_R3 [31:0];
	if(mux_select[4:0] == 5'b00100) BusMuxOut[31:0] <= BusMuxIn_R4 [31:0];
	if(mux_select[4:0] == 5'b00101) BusMuxOut[31:0] <= BusMuxIn_R5 [31:0];
	if(mux_select[4:0] == 5'b00110) BusMuxOut[31:0] <= BusMuxIn_R6 [31:0];
	if(mux_select[4:0] == 5'b00111) BusMuxOut[31:0] <= BusMuxIn_R7 [31:0];
	if(mux_select[4:0] == 5'b01000) BusMuxOut[31:0] <= BusMuxIn_R8 [31:0];
	if(mux_select[4:0] == 5'b01001) BusMuxOut[31:0] <= BusMuxIn_R9 [31:0];
	if(mux_select[4:0] == 5'b01010) BusMuxOut[31:0] <= BusMuxIn_R10 [31:0];
	if(mux_select[4:0] == 5'b01011) BusMuxOut[31:0] <= BusMuxIn_R11 [31:0];
	if(mux_select[4:0] == 5'b01100) BusMuxOut[31:0] <= BusMuxIn_R12 [31:0];
	if(mux_select[4:0] == 5'b01101) BusMuxOut[31:0] <= BusMuxIn_R13 [31:0];
	if(mux_select[4:0] == 5'b01110) BusMuxOut[31:0] <= BusMuxIn_R14 [31:0];
	if(mux_select[4:0] == 5'b01111) BusMuxOut[31:0] <= BusMuxIn_R15 [31:0];
	if(mux_select[4:0] == 5'b10000) BusMuxOut[31:0] <= BusMuxIn_HI [31:0];
	if(mux_select[4:0] == 5'b10001) BusMuxOut[31:0] <= BuxMuxIn_LO [31:0];
	if(mux_select[4:0] == 5'b10010) BusMuxOut[31:0] <= BuxMuxIn_Zhigh [31:0];
	if(mux_select[4:0] == 5'b10011) BusMuxOut[31:0] <= BuxMuxIn_Zlow [31:0];
	if(mux_select[4:0] == 5'b10100) BusMuxOut[31:0] <= BuxMuxIn_PC [31:0];
	if(mux_select[4:0] == 5'b10101) BusMuxOut[31:0] <= BuxMuxIn_MDR [31:0];
	if(mux_select[4:0] == 5'b10110) BusMuxOut[31:0] <= BuxMuxIn_InPort [31:0];
	if(mux_select[4:0] == 5'b10111) BusMuxOut[31:0] <= C_sign_extended [31:0];
	// bit value 24+ unused
	if(mux_select[4:0] == 5'b11000) BusMuxOut[31:0] <= 32'h0;	
	if(mux_select[4:0] == 5'b11001) BusMuxOut[31:0] <= 32'h0;	
	if(mux_select[4:0] == 5'b11010) BusMuxOut[31:0] <= 32'h0;	
	if(mux_select[4:0] == 5'b11011) BusMuxOut[31:0] <= 32'h0;	
	if(mux_select[4:0] == 5'b11100) BusMuxOut[31:0] <= 32'h0;	
	if(mux_select[4:0] == 5'b11101) BusMuxOut[31:0] <= 32'h0;	
	if(mux_select[4:0] == 5'b11110) BusMuxOut[31:0] <= 32'h0;	
	if(mux_select[4:0] == 5'b11111) BusMuxOut[31:0] <= 32'h0;	
end
endmodule