library verilog;
use verilog.vl_types.all;
entity enc_32_to_1_tb is
end enc_32_to_1_tb;
