`timescale 1ns / 10ps
module alu_add(
	input wire[31:0] A,
	input wire [31:0] B,
	output reg [31:0] C
);



endmodule