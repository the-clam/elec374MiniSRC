module seven_seg_out(
    output reg [7:0] display,
    input wire clk,
    input wire [3:0] data
);

always@(negedge clk)
begin
    case(data[3:0])
        4'b0000 : display <= 8'b11000000;
        4'b0001 : display <= 8'b11111001;
        4'b0010 : display <= 8'b10100100;
        4'b0011 : display <= 8'b10110000;
        4'b0100 : display <= 8'b10011001;
        4'b0101 : display <= 8'b10010010;
        4'b0110 : display <= 8'b10000010;
        4'b0111 : display <= 8'b11111000;
        4'b1000 : display <= 8'b10000000;
        4'b1001 : display <= 8'b10010000;
        4'b1010 : display <= 8'b10001000;
        4'b1011 : display <= 8'b10000011;
        4'b1100 : display <= 8'b11000110;
        4'b1101 : display <= 8'b10100001;
        4'b1110 : display <= 8'b10000110;
        4'b1111 : display <= 8'b10001110;
    endcase
end
endmodule
