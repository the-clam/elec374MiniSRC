module dec_4_to_16(
    input wire [3:0] dec_input,
    output reg [15:0] dec_output
);
    always@(*)
    begin
        case(dec_input)
            4'b0000 : dec_output = 16'b0000000000000001;
            4'b0001 : dec_output = 16'b0000000000000010;
            4'b0010 : dec_output = 16'b0000000000000100;
            4'b0011 : dec_output = 16'b0000000000001000;
            4'b0100 : dec_output = 16'b0000000000010000;
            4'b0101 : dec_output = 16'b0000000000100000;
            4'b0110 : dec_output = 16'b0000000001000000;
            4'b0111 : dec_output = 16'b0000000010000000;
            4'b1000 : dec_output = 16'b0000000100000000;
            4'b1001 : dec_output = 16'b0000001000000000;
            4'b1010 : dec_output = 16'b0000010000000000;
            4'b1011 : dec_output = 16'b0000100000000000;
            4'b1100 : dec_output = 16'b0001000000000000;
            4'b1101 : dec_output = 16'b0010000000000000;
            4'b1110 : dec_output = 16'b0100000000000000;
            4'b1111 : dec_output = 16'b1000000000000000;
        endcase
    end
endmodule