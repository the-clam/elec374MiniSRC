`timescale 1ns / 10ps
module alu_mul(
	input wire [31:0] A, // multiplicand
   input wire [31:0] B, // multiplier
	output wire [63:0] P
);

endmodule
