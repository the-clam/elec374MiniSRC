library verilog;
use verilog.vl_types.all;
entity enc_32_to_1 is
    port(
        mux_input_0     : in     vl_logic_vector(31 downto 0);
        mux_input_1     : in     vl_logic_vector(31 downto 0);
        mux_input_2     : in     vl_logic_vector(31 downto 0);
        mux_input_3     : in     vl_logic_vector(31 downto 0);
        mux_input_4     : in     vl_logic_vector(31 downto 0);
        mux_input_5     : in     vl_logic_vector(31 downto 0);
        mux_input_6     : in     vl_logic_vector(31 downto 0);
        mux_input_7     : in     vl_logic_vector(31 downto 0);
        mux_input_8     : in     vl_logic_vector(31 downto 0);
        mux_input_9     : in     vl_logic_vector(31 downto 0);
        mux_input_10    : in     vl_logic_vector(31 downto 0);
        mux_input_11    : in     vl_logic_vector(31 downto 0);
        mux_input_12    : in     vl_logic_vector(31 downto 0);
        mux_input_13    : in     vl_logic_vector(31 downto 0);
        mux_input_14    : in     vl_logic_vector(31 downto 0);
        mux_input_15    : in     vl_logic_vector(31 downto 0);
        mux_input_16    : in     vl_logic_vector(31 downto 0);
        mux_input_17    : in     vl_logic_vector(31 downto 0);
        mux_input_18    : in     vl_logic_vector(31 downto 0);
        mux_input_19    : in     vl_logic_vector(31 downto 0);
        mux_input_20    : in     vl_logic_vector(31 downto 0);
        mux_input_21    : in     vl_logic_vector(31 downto 0);
        mux_input_22    : in     vl_logic_vector(31 downto 0);
        mux_input_23    : in     vl_logic_vector(31 downto 0);
        mux_input_24    : in     vl_logic_vector(31 downto 0);
        mux_input_25    : in     vl_logic_vector(31 downto 0);
        mux_input_26    : in     vl_logic_vector(31 downto 0);
        mux_input_27    : in     vl_logic_vector(31 downto 0);
        mux_input_28    : in     vl_logic_vector(31 downto 0);
        mux_input_29    : in     vl_logic_vector(31 downto 0);
        mux_input_30    : in     vl_logic_vector(31 downto 0);
        mux_input_31    : in     vl_logic_vector(31 downto 0);
        mux_sel         : in     vl_logic_vector(4 downto 0);
        mux_out         : out    vl_logic_vector(31 downto 0)
    );
end enc_32_to_1;
