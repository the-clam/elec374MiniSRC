library verilog;
use verilog.vl_types.all;
entity reg32_tb is
end reg32_tb;
