`timescale 1ns / 10 ps
module alu_add (

);